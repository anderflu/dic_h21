// Module for the 2 x 2 pixel array using pixelSensor

module pixelArray;


    logic [7:0] pixArr [0:1][0:1];






endmodule
